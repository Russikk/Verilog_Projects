`timescale 1ns/1ns

module regFile_tb;

  reg           i_clk, i_we;
  reg   [4:0]   i_raddr1, i_raddr2, i_waddr;
  reg   [31:0]  i_wdata;           
  wire  [31:0]  o_rdata1, o_rdata2;


reg [31:0] registers [31:0];
reg          write_occurred; 

  regFile uut (
    .i_clk(i_clk),
    .i_we(i_we),
    .i_raddr1(i_raddr1),
    .i_raddr2(i_raddr2),
    .i_waddr(i_waddr),
    .i_wdata(i_wdata),
    .o_rdata1(o_rdata1),
    .o_rdata2(o_rdata2)
  );

  // ???????? ?????? ? ???????? 10 ??
  always #5 i_clk = ~i_clk;

  initial begin
    // ????????? ????????
    i_clk = 0;
    i_we = 0;
    i_raddr1 = 5'b0;
    i_raddr2 = 5'b0;
    i_waddr = 5'b0;
    i_wdata = 32'h0000_0000;

    // ????????? ???? ? ???????
    i_waddr = 5'd5;
    i_wdata = 32'h1234_5678;
    i_we = 1;
    #10;
   

    // ???????? ???? ???? ??? ???????? ????
    #10;

    // ??????? ???? ? ????????
    i_raddr1 = 5'd5;
    #10;
  
    i_raddr2 = 5'd0;
    #10;

    // ?????????? ?????????
    $finish;
  end

endmodule

